module logic_andx (input a, b, output out);
 assign out = a & b;
endmodule

module andx (input vd978da, vf5c2a1, output v2a11a2);
 wire w0;
 wire w1;
 wire w2;
 assign w0 = vd978da;
 assign w1 = vf5c2a1;
 assign v2a11a2 = w2;
 logic_andx vf8c369 (
   .a(w0),
   .b(w1),
   .out(w2)
 );
endmodule
