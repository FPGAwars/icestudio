// Generated verilog

module driver0x(output o0);
assign o0 = 1'b0;
endmodule

module main(output output17);
wire w0;
assign output17 = w0;
driver0x driver022 (
    .o0(w0)
);
endmodule
