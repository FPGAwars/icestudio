// Generated verilog

module driver1x(output o0);
assign o0 = 1'b1;
endmodule

module main(output output11);
wire w0;
assign output11 = w0;
driver1x driver110 (
    .o0(w0)
);
endmodule
