// Generated verilog

module main();
endmodule
