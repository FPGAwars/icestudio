module main_vf83e2f (input a, output c);
 // NOT logic gate
 assign c = ! a;
endmodule

module main (input v6c94be, output v3d2176);
 wire w0;
 wire w1;
 assign w0 = v6c94be;
 assign v3d2176 = w1;
 main_vf83e2f v158fc7 (
   .a(w0),
   .c(w1)
 );
endmodule
