module orx (input a, b, output o);
assign o = a | b;
endmodule
