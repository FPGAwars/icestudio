module main_v325b6b_vf83e2f (output v);
 // Driver low
 assign v = 1'b0;
endmodule

module main_v325b6b (output vec9ea9);
 wire w0;
 assign vec9ea9 = w0;
 main_v325b6b_vf83e2f vf9452a (
   .v(w0)
 );
endmodule

module main (output va7d04c);
 wire w0;
 assign va7d04c = w0;
 main_v325b6b vb59771 (
   .vec9ea9(w0)
 );
endmodule
