module driver_driver1x (output out);
 assign out = 1'b1;
endmodule

module highx (output vce929a);
 wire w0;
 assign vce929a = w0;
 driver_driver1x vdfd4f7 (
   .out(w0)
 );
endmodule
