module main (input v0e28cb,
             output vcbab45);
 wire w0;
 wire w1;
 assign w0 = v0e28cb;
 assign vcbab45 = w1;
 main_basic_code_vd54ca1 vd54ca1 (
  .a(w0),
  .c(w1)
 );
endmodule

module main_basic_code_vd54ca1 (input a,
                                output c);
 // NOT logic gate
 
 assign c = ! a;
endmodule

