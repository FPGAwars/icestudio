module vf9452a (output v);
 // Driver low
 assign v = 1'b0;
endmodule

module vb59771 (output vec9ea9);
 wire w0;
 assign vec9ea9 = w0;
 vf9452a vf9452a (
   .v(w0)
 );
endmodule

module main (output va7d04c);
 wire w0;
 assign va7d04c = w0;
 vb59771 vb59771 (
   .vec9ea9(w0)
 );
endmodule
