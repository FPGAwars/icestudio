module driver #(parameter B = 1'b0)(output o);
assign o = B;
endmodule
