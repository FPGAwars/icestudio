module notx (input i, output o);
assign o = ! i;
endmodule
