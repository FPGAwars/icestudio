module main_vf83e2f (input a, input b, output c);
 // OR logic gate
 assign c = a | b;
endmodule

module main (input v0e28cb, input v3ca442, output vcbab45);
 wire w0;
 wire w1;
 wire w2;
 assign w0 = v0e28cb;
 assign w1 = v3ca442;
 assign vcbab45 = w2;
 main_vf83e2f vf4938a (
   .a(w0),
   .b(w1),
   .c(w2)
 );
endmodule
